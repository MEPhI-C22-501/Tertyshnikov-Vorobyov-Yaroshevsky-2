library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package inst_mem_pkg is
    type memory_array is array (0 to 65535) of std_logic_vector(31 downto 0);
end inst_mem_pkg;

package body inst_mem_pkg is
end inst_mem_pkg;
