library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package register_file_pkg is
    type registers_array is array (31 downto 0) of std_logic_vector(31 downto 0);
end register_file_pkg;

package body register_file_pkg is
end register_file_pkg;
