library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package csr_mem_pkg is
    type csr_array is array (31 downto 0) of std_logic_vector(31 downto 0);
end csr_mem_pkg;

package body csr_mem_pkg is
end csr_mem_pkg;
